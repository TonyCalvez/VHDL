library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bascule_d_tb is
end entity;

architecture bhv of bascule_d_tb is

  constant HALF_PERIOD : time := 5 ns;
  signal reset_n : std_logic := '0';
  signal sreset  : std_logic := '0';
  signal running : boolean   := true;

  signal clk    : std_logic := '0';
  signal input  : std_logic := '1';
  signal output : std_logic := '0';
  
  procedure wait_cycles(n : natural) is
   begin
     for i in 1 to n loop
       wait until rising_edge(clk);
     end loop;
   end procedure;



begin
  -------------------------------------------------------------------
  -- clock and reset
  -------------------------------------------------------------------
  reset_n <= '0','1' after 666 ns;
  clk <= not(clk) after HALF_PERIOD when running else clk;

  --------------------------------------------------------------------
  -- Design Under Test
  --------------------------------------------------------------------
  dut : entity work.bascule_d(using_rising_edge)
        
        port map (
          clk    => clk   ,
          input  => input ,
          output => output
        );

  --------------------------------------------------------------------
  -- sequential stimuli
  --------------------------------------------------------------------
  stim : process
   begin
     report "running testbench for bascule_d(using_rising_edge)";
     report "waiting for asynchronous reset";
     wait until reset_n='1';
     wait_cycles(100);
     report "end of simulation";
     running <=false;
     wait;
   end process;

end bhv;
