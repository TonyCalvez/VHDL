library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity counter_enable_tb is
end entity;

architecture bhv of counter_enable_tb is

  constant HALF_PERIOD : time := 5 ns;
  
  signal clk     : std_logic := '0';
  signal reset_n : std_logic := '0';
  signal sreset  : std_logic := '0';
  signal running : boolean   := true;

  procedure wait_cycles(n : natural) is
   begin
     for i in 1 to n loop
       wait until rising_edge(clk);
     end loop;
   end procedure;

  signal enable  : std_logic := '0';
  signal msb     : std_logic := '0';

begin
  -------------------------------------------------------------------
  -- clock and reset
  -------------------------------------------------------------------
  reset_n <= '0','1' after 666 ns;
  enable <= '0','1' after 700 ns;
  clk <= not(clk) after HALF_PERIOD when running else clk;

  --------------------------------------------------------------------
  -- Design Under Test
  --------------------------------------------------------------------
  dut : entity work.counter_enable(rtl)
        port map (
          reset_n => reset_n,
          clk     => clk    ,
          enable  => enable ,
          msb     => msb    
        );

  --------------------------------------------------------------------
  -- sequential stimuli
  --------------------------------------------------------------------
  stim : process
   begin
     report "running testbench for counter_enable(rtl)";
     report "waiting for asynchronous reset";
     wait until reset_n='1';
     wait_cycles(100);
     report "applying stimuli...";
     wait_cycles(100);
     report "end of simulation";
     running <=false;
     wait;
   end process;

end bhv;
